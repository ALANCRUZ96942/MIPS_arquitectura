-------------------------------------------------------------------------------
--
-- Title       : instructionmemory
-- Design      : instructionmemory
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\instructionmemory\instructionmemory\src\instructionmemory.vhd
-- Generated   : Mon Apr 18 23:38:52 2022
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {instructionmemory} architecture {instructionmemory}}

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity InstructionMemory is
	 Generic (size: integer := 32);
    Port (
		AddressIM : in  STD_LOGIC_VECTOR(size-1 downto 0);
		Instruction : out STD_LOGIC_VECTOR (size-1 downto 0);
		Clock : in STD_LOGIC);
end InstructionMemory;

architecture Behavioral of InstructionMemory is
type memoryType is array (0 to 63) of STD_LOGIC_VECTOR (31 downto 0);
signal memory : memoryType :=("00000000000000010001000000100000",
"00000000100000110010100000100010",
"00000000110001110100000000100100",
"00000001001010100101100000100101",
"00000001100011010111000000101010",
"00000001111100001000100000101000",
"10001110010100110000000000000001",
"10101110101101100000000000000001",
"00010000010001010000000000000010",
"10101000000000000000000000000010",
"00000001001000110010100000100000",
"00000000100010010001000000100000",
"00000010000001000010100000100010",
"00000010101100110100000000100100",
"00000001111000010101100000100101",
"00000011111100000111000000101010",
"00000001001000111000100000101000",
"10001100110100110000000000000011",
"10101101111101100000000000000010",
"00010000011100000000000000000101",
"10101000000000000000000000000010",
"00000010000110011000100000100000",
"00000010100111010001000000100000",
"00000010010011110010100000100010",
"00000011000110010100000000100100",
"00000001100011010101100000100101",
"00000010000010100111000000101010",
"00000000011010011000100000101000",
"10001101010100110000000000000100",
"10101111000101100000000000000100",
"00010001100011100000000000000010",
"10101000000000000000000000000100",
"00000001010110110100000000100000",
"00000001111110010001000000100000",
"00000010000001100010100000100010",
"00000000000010010100000000100100",
"00000010100110110101100000100101",
"00000000001000110111000000101010",
"00000011110101011000100000101000",
"10001101010100110000000000000111",
"10101111111101100000000000000111",
"00010000111100000000000000000011",
"10101000000000000000000000000110",
"00000000000111010111000000100000",
"00000001101001100001000000100000",
"00000001101000010010100000100010",
"00000001001111000100000000100100",
"00000001100010010101100000100101",
"00000000100101010111000000101010",
"00000011100010101000100000101000",
"10001110010100110000000000000101",
"10101110111101100000000000000101",
"00010000100000000000000000000111",
"00000010100100000001000000100000",
"00000011001000110010100000100010",
"00000000001001110100000000100100",
"00000011010110110101100000100101",
"00000000000111110111000000101010",
"00000011011111011000100000101000",
"10001100111100110000000000001000",
"10101111110101100000000000001000",
"00010001100100000000000000000100",
"00000011111111010001000000100000",
"00000011001001000010100000100010");
begin
	process(clock)
		begin
			if(rising_edge(clock))then
				if(conv_integer(addressIM(5 downto 0))<64)then
					Instruction <= memory(conv_integer(addressIM(5 downto 0)));
				else
					Instruction <= X"00000000";
				end if;
				--Instruction <= "00000000000000010001000000100000";
			end if;
		end process;
end Behavioral;

